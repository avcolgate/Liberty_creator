VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lib_sample
  CLASS BLOCK ;
  FOREIGN lib_sample ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN BYPASS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.730 11.070 100.000 11.370 ;
    END
  END BYPASS[0]
  PIN BYPASS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.650 77.710 100.000 78.010 ;
    END
  END BYPASS[1]
  PIN BYPASS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.360 82.730 55.500 100.000 ;
    END
  END BYPASS[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.780 0.000 67.920 18.400 ;
    END
  END CLK
  PIN CLK_OUT_DIV
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.590 9.290 88.890 ;
    END
  END CLK_OUT_DIV
  PIN CLK_OUT_G
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.900 86.320 32.040 100.000 ;
    END
  END CLK_OUT_G
  PIN CNTR_OUT1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.160 0.000 0.300 11.600 ;
    END
  END CNTR_OUT1[0]
  PIN CNTR_OUT1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.520 86.320 99.660 100.000 ;
    END
  END CNTR_OUT1[1]
  PIN CNTR_OUT1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.860 0.000 90.000 11.600 ;
    END
  END CNTR_OUT1[2]
  PIN CNTR_OUT2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.240 0.000 22.380 11.600 ;
    END
  END CNTR_OUT2[0]
  PIN CNTR_OUT2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.950 9.290 22.250 ;
    END
  END CNTR_OUT2[1]
  PIN CNTR_OUT2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.990 55.950 100.000 56.250 ;
    END
  END CNTR_OUT2[2]
  PIN CNTR_OUT3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.710 9.290 44.010 ;
    END
  END CNTR_OUT3[0]
  PIN CNTR_OUT3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.440 86.320 77.580 100.000 ;
    END
  END CNTR_OUT3[1]
  PIN CNTR_OUT3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.320 0.000 44.460 11.600 ;
    END
  END CNTR_OUT3[2]
  PIN EN_G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.830 20.790 67.130 ;
    END
  END EN_G
  PIN RST_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.820 76.800 9.960 100.000 ;
    END
  END RST_B
  PIN SELECT_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.270 34.190 100.000 34.490 ;
    END
  END SELECT_3
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.960 10.640 28.560 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.440 10.640 73.040 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.640 94.540 31.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.200 94.540 50.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.760 94.540 70.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.840 10.640 17.440 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.080 10.640 39.680 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.320 10.640 61.920 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.560 10.640 84.160 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.860 94.540 21.460 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 39.420 94.540 41.020 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 58.980 94.540 60.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 78.540 94.540 80.140 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.640 99.750 87.280 ;
      LAYER met2 ;
        RECT 0.100 76.520 9.540 88.925 ;
        RECT 10.240 86.040 31.620 88.925 ;
        RECT 32.320 86.040 55.080 88.925 ;
        RECT 10.240 82.450 55.080 86.040 ;
        RECT 55.780 86.040 77.160 88.925 ;
        RECT 77.860 86.040 99.240 88.925 ;
        RECT 55.780 82.450 99.720 86.040 ;
        RECT 10.240 76.520 99.720 82.450 ;
        RECT 0.100 18.680 99.720 76.520 ;
        RECT 0.100 11.880 67.500 18.680 ;
        RECT 0.580 10.695 21.960 11.880 ;
        RECT 22.660 10.695 44.040 11.880 ;
        RECT 44.740 10.695 67.500 11.880 ;
        RECT 68.200 11.880 99.720 18.680 ;
        RECT 68.200 10.695 89.580 11.880 ;
        RECT 90.280 10.695 99.720 11.880 ;
      LAYER met3 ;
        RECT 9.690 88.190 91.015 88.905 ;
        RECT 9.265 78.410 91.015 88.190 ;
        RECT 9.265 77.310 77.250 78.410 ;
        RECT 9.265 67.530 91.015 77.310 ;
        RECT 21.190 66.430 91.015 67.530 ;
        RECT 9.265 56.650 91.015 66.430 ;
        RECT 9.265 55.550 90.590 56.650 ;
        RECT 9.265 44.410 91.015 55.550 ;
        RECT 9.690 43.310 91.015 44.410 ;
        RECT 9.265 34.890 91.015 43.310 ;
        RECT 9.265 33.790 75.870 34.890 ;
        RECT 9.265 22.650 91.015 33.790 ;
        RECT 9.690 21.550 91.015 22.650 ;
        RECT 9.265 11.770 91.015 21.550 ;
        RECT 9.265 10.715 76.330 11.770 ;
  END
END lib_sample
END LIBRARY

